
LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
 
-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--USE ieee.numeric_std.ALL;
 
ENTITY tb_procesador IS
END tb_procesador;
 
ARCHITECTURE behavior OF tb_procesador IS 
 
    -- Component Declaration for the Unit Under Test (UUT)

    COMPONENT primerprocesador
    PORT(
         clk : IN  std_logic;
         rst : IN  std_logic;
         resultado : OUT  std_logic_vector(31 downto 0)
        );
    END COMPONENT;
    

   --Inputs
   signal clk : std_logic := '0';
   signal rst : std_logic := '0';

 	--Outputs
   signal resultado : std_logic_vector(31 downto 0);

   -- Clock period definitions
   constant clk_period : time := 10 ns;
 
BEGIN
 
	-- Instantiate the Unit Under Test (UUT)
   uut: primerprocesador PORT MAP (
          clk => clk,
          rst => rst,
          resultado => resultado
        );

   -- Clock process definitions
   clk_process :process
   begin



		clk <= '0';
		wait for clk_period/2;
		clk <= '1';
		wait for clk_period/2;
   end process;
 

   -- Stimulus process
   stim_proc: process
   begin		
		wait for 10 ns;
      rst <= '1';
      wait for 10 ns;	
		rst <= '0';
      wait;
   end process;

END;
